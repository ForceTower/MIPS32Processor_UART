module Processador(input clock);
	reg [31:0] pc;
	initial begin
		pc <= 32'd0;
	end
endmodule 